library ieee;
use ieee.std_logic_1164.all; 
use ieee.std_logic_unsigned.all;

entity ROM_176x4 is
  port (Clock : in std_logic;
  		CS_L : in std_logic;
        R_W  : in std_logic;
        Addr   : in std_logic_vector(7 downto 0);
        Data  : out std_logic_vector(3 downto 0));
end ROM_176x4;

architecture ROM_176x4_Arch of ROM_176x4 is
  type rom_type is array (0 to 175)
        of std_logic_vector (3 downto 0);
  signal ROM : rom_type;
  signal Read_Enable : std_logic;
begin

ROM(0) <= X"7";
ROM(1) <= X"0";
ROM(2) <= X"D";
ROM(3) <= X"0";
ROM(4) <= X"B";
ROM(5) <= X"7";
ROM(6) <= X"1";
ROM(7) <= X"D";
ROM(8) <= X"1";
ROM(9) <= X"B";
ROM(10) <= X"9";
ROM(11) <= X"D";
ROM(12) <= X"5";
ROM(13) <= X"F";
ROM(14) <= X"1";
ROM(15) <= X"B";
ROM(16) <= X"6";
ROM(17) <= X"7";
ROM(18) <= X"A";
ROM(19) <= X"D";
ROM(20) <= X"1";
ROM(21) <= X"6";
ROM(22) <= X"A";
ROM(23) <= X"D";
ROM(24) <= X"1";
ROM(25) <= X"B";
ROM(26) <= X"9";
ROM(27) <= X"2";
ROM(28) <= X"2";
ROM(29) <= X"7";
ROM(30) <= X"1";
ROM(31) <= X"D";
ROM(32) <= X"1";
ROM(33) <= X"B";
ROM(34) <= X"5";
ROM(35) <= X"0";
ROM(36) <= X"6";
ROM(37) <= X"F";
ROM(38) <= X"A";
ROM(39) <= X"3";
ROM(40) <= X"3";
ROM(41) <= X"5";
ROM(42) <= X"1";
ROM(43) <= X"6";
ROM(44) <= X"F";
ROM(45) <= X"A";
ROM(46) <= X"3";
ROM(47) <= X"3";
ROM(48) <= X"9";
ROM(49) <= X"D";
ROM(50) <= X"5";
ROM(51) <= X"5";
ROM(52) <= X"0";
ROM(53) <= X"A";
ROM(54) <= X"0";
ROM(55) <= X"4";
ROM(56) <= X"5";
ROM(57) <= X"1";
ROM(58) <= X"A";
ROM(59) <= X"D";
ROM(60) <= X"4";
ROM(61) <= X"9";
ROM(62) <= X"D";
ROM(63) <= X"5";
ROM(64) <= X"F";
ROM(65) <= X"0";
ROM(66) <= X"B";
ROM(67) <= X"6";
ROM(68) <= X"D";
ROM(69) <= X"A";
ROM(70) <= X"A";
ROM(71) <= X"5";
ROM(72) <= X"6";
ROM(73) <= X"4";
ROM(74) <= X"9";
ROM(75) <= X"A";
ROM(76) <= X"5";
ROM(77) <= X"F";
ROM(78) <= X"0";
ROM(79) <= X"B";
ROM(80) <= X"A";
ROM(81) <= X"8";
ROM(82) <= X"5";
ROM(83) <= X"6";
ROM(84) <= X"F";
ROM(85) <= X"9";
ROM(86) <= X"A";
ROM(87) <= X"5";
ROM(88) <= X"7";
ROM(89) <= X"3";
ROM(90) <= X"D";
ROM(91) <= X"0";
ROM(92) <= X"B";
ROM(93) <= X"F";
ROM(94) <= X"0";
ROM(95) <= X"B";
ROM(96) <= X"A";
ROM(97) <= X"6";
ROM(98) <= X"9";
ROM(99) <= X"6";
ROM(100) <= X"F";
ROM(101) <= X"A";
ROM(102) <= X"A";
ROM(103) <= X"8";
ROM(104) <= X"6";
ROM(105) <= X"F";
ROM(106) <= X"A";
ROM(107) <= X"E";
ROM(108) <= X"7";
ROM(109) <= X"6";
ROM(110) <= X"F";
ROM(111) <= X"A";
ROM(112) <= X"2";
ROM(113) <= X"7";
ROM(114) <= X"4";
ROM(115) <= X"0";
ROM(116) <= X"4";
ROM(117) <= X"2";
ROM(118) <= X"F";
ROM(119) <= X"1";
ROM(120) <= X"B";
ROM(121) <= X"4";
ROM(122) <= X"3";
ROM(123) <= X"9";
ROM(124) <= X"D";
ROM(125) <= X"0";
ROM(126) <= X"4";
ROM(127) <= X"1";
ROM(128) <= X"4";
ROM(129) <= X"3";
ROM(130) <= X"F";
ROM(131) <= X"1";
ROM(132) <= X"B";
ROM(133) <= X"4";
ROM(134) <= X"2";
ROM(135) <= X"9";
ROM(136) <= X"D";
ROM(137) <= X"0";
ROM(138) <= X"4";
ROM(139) <= X"0";
ROM(140) <= X"4";
ROM(141) <= X"2";
ROM(142) <= X"F";
ROM(143) <= X"1";
ROM(144) <= X"B";
ROM(145) <= X"4";
ROM(146) <= X"1";
ROM(147) <= X"9";
ROM(148) <= X"D";
ROM(149) <= X"0";
ROM(150) <= X"4";
ROM(151) <= X"1";
ROM(152) <= X"4";
ROM(153) <= X"3";
ROM(154) <= X"F";
ROM(155) <= X"1";
ROM(156) <= X"B";
ROM(157) <= X"4";
ROM(158) <= X"0";
ROM(159) <= X"9";
ROM(160) <= X"D";
ROM(161) <= X"0";
ROM(162) <= X"0";
ROM(163) <= X"0";
ROM(164) <= X"0";
ROM(165) <= X"0";
ROM(166) <= X"0";
ROM(167) <= X"0";
ROM(168) <= X"0";
ROM(169) <= X"0";
ROM(170) <= X"0";
ROM(171) <= X"0";
ROM(172) <= X"0";
ROM(173) <= X"0";
ROM(174) <= X"0";
ROM(175) <= X"0";
	Read_Enable <=  '0' when(CS_L='0' and R_W = '1') else '1';

	process (Clock)
	begin
		if(Clock='0') then
			if(Read_Enable = '0') then
			  Data  <= ROM(conv_integer(Addr));
		  	else
			  Data <= "ZZZZ";
	      	end if;
		else Data <= "ZZZZ";
		end if;

	end process;

	end ROM_176x4_Arch;
